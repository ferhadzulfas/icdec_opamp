magic
tech sky130A
magscale 1 2
timestamp 1729236971
<< error_p >>
rect -988 181 -916 187
rect -716 181 -644 187
rect -444 181 -372 187
rect -172 181 -100 187
rect 100 181 172 187
rect 372 181 444 187
rect 644 181 716 187
rect 916 181 988 187
rect -988 147 -976 181
rect -716 147 -704 181
rect -444 147 -432 181
rect -172 147 -160 181
rect 100 147 112 181
rect 372 147 384 181
rect 644 147 656 181
rect 916 147 928 181
rect -988 141 -916 147
rect -716 141 -644 147
rect -444 141 -372 147
rect -172 141 -100 147
rect 100 141 172 147
rect 372 141 444 147
rect 644 141 716 147
rect 916 141 988 147
rect -988 -147 -916 -141
rect -716 -147 -644 -141
rect -444 -147 -372 -141
rect -172 -147 -100 -141
rect 100 -147 172 -141
rect 372 -147 444 -141
rect 644 -147 716 -141
rect 916 -147 988 -141
rect -988 -181 -976 -147
rect -716 -181 -704 -147
rect -444 -181 -432 -147
rect -172 -181 -160 -147
rect 100 -181 112 -147
rect 372 -181 384 -147
rect 644 -181 656 -147
rect 916 -181 928 -147
rect -988 -187 -916 -181
rect -716 -187 -644 -181
rect -444 -187 -372 -181
rect -172 -187 -100 -181
rect 100 -187 172 -181
rect 372 -187 444 -181
rect 644 -187 716 -181
rect 916 -187 988 -181
<< nwell >>
rect -1096 -200 1096 200
<< pmos >>
rect -1002 -100 -902 100
rect -730 -100 -630 100
rect -458 -100 -358 100
rect -186 -100 -86 100
rect 86 -100 186 100
rect 358 -100 458 100
rect 630 -100 730 100
rect 902 -100 1002 100
<< pdiff >>
rect -1060 88 -1002 100
rect -1060 -88 -1048 88
rect -1014 -88 -1002 88
rect -1060 -100 -1002 -88
rect -902 88 -844 100
rect -902 -88 -890 88
rect -856 -88 -844 88
rect -902 -100 -844 -88
rect -788 88 -730 100
rect -788 -88 -776 88
rect -742 -88 -730 88
rect -788 -100 -730 -88
rect -630 88 -572 100
rect -630 -88 -618 88
rect -584 -88 -572 88
rect -630 -100 -572 -88
rect -516 88 -458 100
rect -516 -88 -504 88
rect -470 -88 -458 88
rect -516 -100 -458 -88
rect -358 88 -300 100
rect -358 -88 -346 88
rect -312 -88 -300 88
rect -358 -100 -300 -88
rect -244 88 -186 100
rect -244 -88 -232 88
rect -198 -88 -186 88
rect -244 -100 -186 -88
rect -86 88 -28 100
rect -86 -88 -74 88
rect -40 -88 -28 88
rect -86 -100 -28 -88
rect 28 88 86 100
rect 28 -88 40 88
rect 74 -88 86 88
rect 28 -100 86 -88
rect 186 88 244 100
rect 186 -88 198 88
rect 232 -88 244 88
rect 186 -100 244 -88
rect 300 88 358 100
rect 300 -88 312 88
rect 346 -88 358 88
rect 300 -100 358 -88
rect 458 88 516 100
rect 458 -88 470 88
rect 504 -88 516 88
rect 458 -100 516 -88
rect 572 88 630 100
rect 572 -88 584 88
rect 618 -88 630 88
rect 572 -100 630 -88
rect 730 88 788 100
rect 730 -88 742 88
rect 776 -88 788 88
rect 730 -100 788 -88
rect 844 88 902 100
rect 844 -88 856 88
rect 890 -88 902 88
rect 844 -100 902 -88
rect 1002 88 1060 100
rect 1002 -88 1014 88
rect 1048 -88 1060 88
rect 1002 -100 1060 -88
<< pdiffc >>
rect -1048 -88 -1014 88
rect -890 -88 -856 88
rect -776 -88 -742 88
rect -618 -88 -584 88
rect -504 -88 -470 88
rect -346 -88 -312 88
rect -232 -88 -198 88
rect -74 -88 -40 88
rect 40 -88 74 88
rect 198 -88 232 88
rect 312 -88 346 88
rect 470 -88 504 88
rect 584 -88 618 88
rect 742 -88 776 88
rect 856 -88 890 88
rect 1014 -88 1048 88
<< poly >>
rect -1002 181 -902 197
rect -1002 147 -986 181
rect -918 147 -902 181
rect -1002 100 -902 147
rect -730 181 -630 197
rect -730 147 -714 181
rect -646 147 -630 181
rect -730 100 -630 147
rect -458 181 -358 197
rect -458 147 -442 181
rect -374 147 -358 181
rect -458 100 -358 147
rect -186 181 -86 197
rect -186 147 -170 181
rect -102 147 -86 181
rect -186 100 -86 147
rect 86 181 186 197
rect 86 147 102 181
rect 170 147 186 181
rect 86 100 186 147
rect 358 181 458 197
rect 358 147 374 181
rect 442 147 458 181
rect 358 100 458 147
rect 630 181 730 197
rect 630 147 646 181
rect 714 147 730 181
rect 630 100 730 147
rect 902 181 1002 197
rect 902 147 918 181
rect 986 147 1002 181
rect 902 100 1002 147
rect -1002 -147 -902 -100
rect -1002 -181 -986 -147
rect -918 -181 -902 -147
rect -1002 -197 -902 -181
rect -730 -147 -630 -100
rect -730 -181 -714 -147
rect -646 -181 -630 -147
rect -730 -197 -630 -181
rect -458 -147 -358 -100
rect -458 -181 -442 -147
rect -374 -181 -358 -147
rect -458 -197 -358 -181
rect -186 -147 -86 -100
rect -186 -181 -170 -147
rect -102 -181 -86 -147
rect -186 -197 -86 -181
rect 86 -147 186 -100
rect 86 -181 102 -147
rect 170 -181 186 -147
rect 86 -197 186 -181
rect 358 -147 458 -100
rect 358 -181 374 -147
rect 442 -181 458 -147
rect 358 -197 458 -181
rect 630 -147 730 -100
rect 630 -181 646 -147
rect 714 -181 730 -147
rect 630 -197 730 -181
rect 902 -147 1002 -100
rect 902 -181 918 -147
rect 986 -181 1002 -147
rect 902 -197 1002 -181
<< polycont >>
rect -986 147 -918 181
rect -714 147 -646 181
rect -442 147 -374 181
rect -170 147 -102 181
rect 102 147 170 181
rect 374 147 442 181
rect 646 147 714 181
rect 918 147 986 181
rect -986 -181 -918 -147
rect -714 -181 -646 -147
rect -442 -181 -374 -147
rect -170 -181 -102 -147
rect 102 -181 170 -147
rect 374 -181 442 -147
rect 646 -181 714 -147
rect 918 -181 986 -147
<< locali >>
rect -1002 147 -986 181
rect -918 147 -902 181
rect -730 147 -714 181
rect -646 147 -630 181
rect -458 147 -442 181
rect -374 147 -358 181
rect -186 147 -170 181
rect -102 147 -86 181
rect 86 147 102 181
rect 170 147 186 181
rect 358 147 374 181
rect 442 147 458 181
rect 630 147 646 181
rect 714 147 730 181
rect 902 147 918 181
rect 986 147 1002 181
rect -1048 88 -1014 104
rect -1048 -104 -1014 -88
rect -890 88 -856 104
rect -890 -104 -856 -88
rect -776 88 -742 104
rect -776 -104 -742 -88
rect -618 88 -584 104
rect -618 -104 -584 -88
rect -504 88 -470 104
rect -504 -104 -470 -88
rect -346 88 -312 104
rect -346 -104 -312 -88
rect -232 88 -198 104
rect -232 -104 -198 -88
rect -74 88 -40 104
rect -74 -104 -40 -88
rect 40 88 74 104
rect 40 -104 74 -88
rect 198 88 232 104
rect 198 -104 232 -88
rect 312 88 346 104
rect 312 -104 346 -88
rect 470 88 504 104
rect 470 -104 504 -88
rect 584 88 618 104
rect 584 -104 618 -88
rect 742 88 776 104
rect 742 -104 776 -88
rect 856 88 890 104
rect 856 -104 890 -88
rect 1014 88 1048 104
rect 1014 -104 1048 -88
rect -1002 -181 -986 -147
rect -918 -181 -902 -147
rect -730 -181 -714 -147
rect -646 -181 -630 -147
rect -458 -181 -442 -147
rect -374 -181 -358 -147
rect -186 -181 -170 -147
rect -102 -181 -86 -147
rect 86 -181 102 -147
rect 170 -181 186 -147
rect 358 -181 374 -147
rect 442 -181 458 -147
rect 630 -181 646 -147
rect 714 -181 730 -147
rect 902 -181 918 -147
rect 986 -181 1002 -147
<< viali >>
rect -976 147 -928 181
rect -704 147 -656 181
rect -432 147 -384 181
rect -160 147 -112 181
rect 112 147 160 181
rect 384 147 432 181
rect 656 147 704 181
rect 928 147 976 181
rect -1048 -88 -1014 88
rect -890 -88 -856 88
rect -776 -88 -742 88
rect -618 -88 -584 88
rect -504 -88 -470 88
rect -346 -88 -312 88
rect -232 -88 -198 88
rect -74 -88 -40 88
rect 40 -88 74 88
rect 198 -88 232 88
rect 312 -88 346 88
rect 470 -88 504 88
rect 584 -88 618 88
rect 742 -88 776 88
rect 856 -88 890 88
rect 1014 -88 1048 88
rect -976 -181 -928 -147
rect -704 -181 -656 -147
rect -432 -181 -384 -147
rect -160 -181 -112 -147
rect 112 -181 160 -147
rect 384 -181 432 -147
rect 656 -181 704 -147
rect 928 -181 976 -147
<< metal1 >>
rect -988 181 -916 187
rect -988 147 -976 181
rect -928 147 -916 181
rect -988 141 -916 147
rect -716 181 -644 187
rect -716 147 -704 181
rect -656 147 -644 181
rect -716 141 -644 147
rect -444 181 -372 187
rect -444 147 -432 181
rect -384 147 -372 181
rect -444 141 -372 147
rect -172 181 -100 187
rect -172 147 -160 181
rect -112 147 -100 181
rect -172 141 -100 147
rect 100 181 172 187
rect 100 147 112 181
rect 160 147 172 181
rect 100 141 172 147
rect 372 181 444 187
rect 372 147 384 181
rect 432 147 444 181
rect 372 141 444 147
rect 644 181 716 187
rect 644 147 656 181
rect 704 147 716 181
rect 644 141 716 147
rect 916 181 988 187
rect 916 147 928 181
rect 976 147 988 181
rect 916 141 988 147
rect -1054 88 -1008 100
rect -1054 -88 -1048 88
rect -1014 -88 -1008 88
rect -1054 -100 -1008 -88
rect -896 88 -850 100
rect -896 -88 -890 88
rect -856 -88 -850 88
rect -896 -100 -850 -88
rect -782 88 -736 100
rect -782 -88 -776 88
rect -742 -88 -736 88
rect -782 -100 -736 -88
rect -624 88 -578 100
rect -624 -88 -618 88
rect -584 -88 -578 88
rect -624 -100 -578 -88
rect -510 88 -464 100
rect -510 -88 -504 88
rect -470 -88 -464 88
rect -510 -100 -464 -88
rect -352 88 -306 100
rect -352 -88 -346 88
rect -312 -88 -306 88
rect -352 -100 -306 -88
rect -238 88 -192 100
rect -238 -88 -232 88
rect -198 -88 -192 88
rect -238 -100 -192 -88
rect -80 88 -34 100
rect -80 -88 -74 88
rect -40 -88 -34 88
rect -80 -100 -34 -88
rect 34 88 80 100
rect 34 -88 40 88
rect 74 -88 80 88
rect 34 -100 80 -88
rect 192 88 238 100
rect 192 -88 198 88
rect 232 -88 238 88
rect 192 -100 238 -88
rect 306 88 352 100
rect 306 -88 312 88
rect 346 -88 352 88
rect 306 -100 352 -88
rect 464 88 510 100
rect 464 -88 470 88
rect 504 -88 510 88
rect 464 -100 510 -88
rect 578 88 624 100
rect 578 -88 584 88
rect 618 -88 624 88
rect 578 -100 624 -88
rect 736 88 782 100
rect 736 -88 742 88
rect 776 -88 782 88
rect 736 -100 782 -88
rect 850 88 896 100
rect 850 -88 856 88
rect 890 -88 896 88
rect 850 -100 896 -88
rect 1008 88 1054 100
rect 1008 -88 1014 88
rect 1048 -88 1054 88
rect 1008 -100 1054 -88
rect -988 -147 -916 -141
rect -988 -181 -976 -147
rect -928 -181 -916 -147
rect -988 -187 -916 -181
rect -716 -147 -644 -141
rect -716 -181 -704 -147
rect -656 -181 -644 -147
rect -716 -187 -644 -181
rect -444 -147 -372 -141
rect -444 -181 -432 -147
rect -384 -181 -372 -147
rect -444 -187 -372 -181
rect -172 -147 -100 -141
rect -172 -181 -160 -147
rect -112 -181 -100 -147
rect -172 -187 -100 -181
rect 100 -147 172 -141
rect 100 -181 112 -147
rect 160 -181 172 -147
rect 100 -187 172 -181
rect 372 -147 444 -141
rect 372 -181 384 -147
rect 432 -181 444 -147
rect 372 -187 444 -181
rect 644 -147 716 -141
rect 644 -181 656 -147
rect 704 -181 716 -147
rect 644 -187 716 -181
rect 916 -147 988 -141
rect 916 -181 928 -147
rect 976 -181 988 -147
rect 916 -187 988 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
