magic
tech sky130A
magscale 1 2
timestamp 1729426932
<< nwell >>
rect -1160 1564 -147 1773
rect 1693 1631 2493 1773
rect 1690 1132 2494 1631
<< viali >>
rect 1339 1378 1579 1618
rect 1339 827 1579 1067
rect 1147 360 1181 481
rect 1341 260 1581 500
rect 1341 -21 1581 219
rect 588 -104 623 -70
<< metal1 >>
rect -331 1698 2075 1732
rect -331 1551 -297 1698
rect 1419 1624 1496 1698
rect 1327 1618 1591 1624
rect 1327 1378 1339 1618
rect 1579 1378 1591 1618
rect 1327 1372 1591 1378
rect 1329 1103 1339 1343
rect 1579 1103 1589 1343
rect 2041 1224 2075 1698
rect 1327 1067 1591 1073
rect -174 976 -164 1041
rect -89 1037 -79 1041
rect -89 992 17 1037
rect -89 976 -79 992
rect -252 890 10 924
rect -252 814 -218 890
rect 1327 827 1339 1067
rect 1579 929 1591 1067
rect 1579 871 1664 929
rect 1579 827 1591 871
rect 1327 821 1591 827
rect -460 768 -318 814
rect -294 768 -218 814
rect 1329 542 1339 782
rect 1579 542 1589 782
rect 1621 526 1663 871
rect 1981 526 2049 567
rect 1329 500 1593 506
rect 1329 493 1341 500
rect 1141 481 1341 493
rect 1141 360 1147 481
rect 1181 360 1341 481
rect 1141 349 1341 360
rect 1141 348 1187 349
rect 588 -64 624 314
rect 1329 260 1341 349
rect 1581 260 1593 500
rect 1621 489 2049 526
rect 1641 391 1651 443
rect 1703 438 1713 443
rect 1703 395 1989 438
rect 1703 391 1713 395
rect 1329 254 1593 260
rect 1329 219 1593 225
rect 1329 -21 1341 219
rect 1581 136 1593 219
rect 1581 75 1704 136
rect 1581 -21 1593 75
rect 1329 -27 1593 -21
rect 576 -70 635 -64
rect 576 -104 588 -70
rect 623 -104 635 -70
rect 576 -110 635 -104
rect 1645 -203 1704 75
rect 1635 -267 1645 -203
rect 1704 -267 1714 -203
<< via1 >>
rect 1339 1103 1579 1343
rect -164 976 -89 1041
rect 1339 542 1579 782
rect 1651 391 1703 443
rect 1645 -267 1704 -203
<< metal2 >>
rect 1339 1343 1579 1353
rect 1245 1278 1287 1279
rect 1245 1226 1339 1278
rect -164 1041 -89 1051
rect 582 992 633 1022
rect 1245 992 1287 1226
rect 1339 1093 1579 1103
rect -164 966 -89 976
rect 581 954 1287 992
rect 582 949 633 954
rect 1339 782 1579 792
rect -946 715 -890 725
rect 1579 596 1663 616
rect 1579 567 1664 596
rect 1339 532 1579 542
rect 1620 453 1664 567
rect 1620 443 1703 453
rect 1620 395 1651 443
rect 1651 381 1703 391
rect -946 329 -890 339
rect 13 95 96 105
rect -430 14 -374 24
rect -331 20 13 92
rect 13 6 96 16
rect 1645 -203 1704 -193
rect 1645 -277 1704 -267
rect -430 -372 -374 -362
rect 1436 -710 1848 -660
<< via2 >>
rect -154 981 -98 1037
rect -946 339 -890 715
rect -430 -362 -374 14
rect 13 16 96 95
rect 1645 -267 1704 -203
<< metal3 >>
rect -164 1037 -88 1042
rect -164 981 -154 1037
rect -98 981 -88 1037
rect -164 976 -88 981
rect -956 715 -880 720
rect -956 339 -946 715
rect -890 339 -880 715
rect -956 334 -880 339
rect -954 204 -881 334
rect -163 204 -93 976
rect -954 144 -93 204
rect -954 142 -364 144
rect -439 19 -364 142
rect -440 14 -364 19
rect -440 -362 -430 14
rect -374 -362 -364 14
rect 3 95 106 100
rect 2065 95 2122 98
rect 3 16 13 95
rect 96 16 2124 95
rect 3 11 106 16
rect 2065 13 2122 16
rect -440 -367 -364 -362
rect 1635 -203 1714 -198
rect 1635 -267 1645 -203
rect 1704 -267 1714 -203
rect 723 -1110 799 -944
rect 1635 -1110 1714 -267
rect 723 -1177 2343 -1110
use nmoscs  nmoscs_0 ~/operationalamplifier/nmoscs
timestamp 1729245215
transform 1 0 205 0 1 365
box -288 -71 976 1265
use nmosdiff  nmosdiff_0 ~/operationalamplifier/nmosdiff
timestamp 1729382277
transform 1 0 131 0 1 -629
box -214 -663 1495 559
use pmoscs  pmoscs_0 ~/operationalamplifier/pmoscs
timestamp 1729158298
transform 1 0 -983 0 1 -1174
box -176 -101 836 2801
use pmosdiff  pmosdiff_0 ~/operationalamplifier/pmosdiff
timestamp 1729387919
transform 1 0 1599 0 1 760
box 94 -2032 894 512
<< labels >>
flabel viali 1479 1485 1479 1485 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel via1 1447 1223 1447 1223 0 FreeSans 1600 0 0 0 RS
port 1 nsew
flabel viali 1463 942 1463 942 0 FreeSans 1600 0 0 0 VIP
port 2 nsew
flabel via1 1465 660 1465 660 0 FreeSans 1600 0 0 0 VIN
port 3 nsew
flabel viali 1468 379 1468 379 0 FreeSans 1600 0 0 0 GND
port 4 nsew
flabel viali 1461 133 1461 133 0 FreeSans 1600 0 0 0 OUT
port 5 nsew
<< end >>
