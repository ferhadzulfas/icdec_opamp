magic
tech sky130A
magscale 1 2
timestamp 1729223494
<< nmos >>
rect -286 727 -86 1127
rect 86 727 286 1127
rect -286 109 -86 509
rect 86 109 286 509
rect -286 -509 -86 -109
rect 86 -509 286 -109
rect -286 -1127 -86 -727
rect 86 -1127 286 -727
<< ndiff >>
rect -344 1115 -286 1127
rect -344 739 -332 1115
rect -298 739 -286 1115
rect -344 727 -286 739
rect -86 1115 -28 1127
rect -86 739 -74 1115
rect -40 739 -28 1115
rect -86 727 -28 739
rect 28 1115 86 1127
rect 28 739 40 1115
rect 74 739 86 1115
rect 28 727 86 739
rect 286 1115 344 1127
rect 286 739 298 1115
rect 332 739 344 1115
rect 286 727 344 739
rect -344 497 -286 509
rect -344 121 -332 497
rect -298 121 -286 497
rect -344 109 -286 121
rect -86 497 -28 509
rect -86 121 -74 497
rect -40 121 -28 497
rect -86 109 -28 121
rect 28 497 86 509
rect 28 121 40 497
rect 74 121 86 497
rect 28 109 86 121
rect 286 497 344 509
rect 286 121 298 497
rect 332 121 344 497
rect 286 109 344 121
rect -344 -121 -286 -109
rect -344 -497 -332 -121
rect -298 -497 -286 -121
rect -344 -509 -286 -497
rect -86 -121 -28 -109
rect -86 -497 -74 -121
rect -40 -497 -28 -121
rect -86 -509 -28 -497
rect 28 -121 86 -109
rect 28 -497 40 -121
rect 74 -497 86 -121
rect 28 -509 86 -497
rect 286 -121 344 -109
rect 286 -497 298 -121
rect 332 -497 344 -121
rect 286 -509 344 -497
rect -344 -739 -286 -727
rect -344 -1115 -332 -739
rect -298 -1115 -286 -739
rect -344 -1127 -286 -1115
rect -86 -739 -28 -727
rect -86 -1115 -74 -739
rect -40 -1115 -28 -739
rect -86 -1127 -28 -1115
rect 28 -739 86 -727
rect 28 -1115 40 -739
rect 74 -1115 86 -739
rect 28 -1127 86 -1115
rect 286 -739 344 -727
rect 286 -1115 298 -739
rect 332 -1115 344 -739
rect 286 -1127 344 -1115
<< ndiffc >>
rect -332 739 -298 1115
rect -74 739 -40 1115
rect 40 739 74 1115
rect 298 739 332 1115
rect -332 121 -298 497
rect -74 121 -40 497
rect 40 121 74 497
rect 298 121 332 497
rect -332 -497 -298 -121
rect -74 -497 -40 -121
rect 40 -497 74 -121
rect 298 -497 332 -121
rect -332 -1115 -298 -739
rect -74 -1115 -40 -739
rect 40 -1115 74 -739
rect 298 -1115 332 -739
<< poly >>
rect -286 1199 -86 1215
rect -286 1165 -270 1199
rect -102 1165 -86 1199
rect -286 1127 -86 1165
rect 86 1199 286 1215
rect 86 1165 102 1199
rect 270 1165 286 1199
rect 86 1127 286 1165
rect -286 689 -86 727
rect -286 655 -270 689
rect -102 655 -86 689
rect -286 639 -86 655
rect 86 689 286 727
rect 86 655 102 689
rect 270 655 286 689
rect 86 639 286 655
rect -286 581 -86 597
rect -286 547 -270 581
rect -102 547 -86 581
rect -286 509 -86 547
rect 86 581 286 597
rect 86 547 102 581
rect 270 547 286 581
rect 86 509 286 547
rect -286 71 -86 109
rect -286 37 -270 71
rect -102 37 -86 71
rect -286 21 -86 37
rect 86 71 286 109
rect 86 37 102 71
rect 270 37 286 71
rect 86 21 286 37
rect -286 -37 -86 -21
rect -286 -71 -270 -37
rect -102 -71 -86 -37
rect -286 -109 -86 -71
rect 86 -37 286 -21
rect 86 -71 102 -37
rect 270 -71 286 -37
rect 86 -109 286 -71
rect -286 -547 -86 -509
rect -286 -581 -270 -547
rect -102 -581 -86 -547
rect -286 -597 -86 -581
rect 86 -547 286 -509
rect 86 -581 102 -547
rect 270 -581 286 -547
rect 86 -597 286 -581
rect -286 -655 -86 -639
rect -286 -689 -270 -655
rect -102 -689 -86 -655
rect -286 -727 -86 -689
rect 86 -655 286 -639
rect 86 -689 102 -655
rect 270 -689 286 -655
rect 86 -727 286 -689
rect -286 -1165 -86 -1127
rect -286 -1199 -270 -1165
rect -102 -1199 -86 -1165
rect -286 -1215 -86 -1199
rect 86 -1165 286 -1127
rect 86 -1199 102 -1165
rect 270 -1199 286 -1165
rect 86 -1215 286 -1199
<< polycont >>
rect -270 1165 -102 1199
rect 102 1165 270 1199
rect -270 655 -102 689
rect 102 655 270 689
rect -270 547 -102 581
rect 102 547 270 581
rect -270 37 -102 71
rect 102 37 270 71
rect -270 -71 -102 -37
rect 102 -71 270 -37
rect -270 -581 -102 -547
rect 102 -581 270 -547
rect -270 -689 -102 -655
rect 102 -689 270 -655
rect -270 -1199 -102 -1165
rect 102 -1199 270 -1165
<< locali >>
rect -286 1165 -270 1199
rect -102 1165 -86 1199
rect 86 1165 102 1199
rect 270 1165 286 1199
rect -332 1115 -298 1131
rect -332 723 -298 739
rect -74 1115 -40 1131
rect -74 723 -40 739
rect 40 1115 74 1131
rect 40 723 74 739
rect 298 1115 332 1131
rect 298 723 332 739
rect -286 655 -270 689
rect -102 655 -86 689
rect 86 655 102 689
rect 270 655 286 689
rect -286 547 -270 581
rect -102 547 -86 581
rect 86 547 102 581
rect 270 547 286 581
rect -332 497 -298 513
rect -332 105 -298 121
rect -74 497 -40 513
rect -74 105 -40 121
rect 40 497 74 513
rect 40 105 74 121
rect 298 497 332 513
rect 298 105 332 121
rect -286 37 -270 71
rect -102 37 -86 71
rect 86 37 102 71
rect 270 37 286 71
rect -286 -71 -270 -37
rect -102 -71 -86 -37
rect 86 -71 102 -37
rect 270 -71 286 -37
rect -332 -121 -298 -105
rect -332 -513 -298 -497
rect -74 -121 -40 -105
rect -74 -513 -40 -497
rect 40 -121 74 -105
rect 40 -513 74 -497
rect 298 -121 332 -105
rect 298 -513 332 -497
rect -286 -581 -270 -547
rect -102 -581 -86 -547
rect 86 -581 102 -547
rect 270 -581 286 -547
rect -286 -689 -270 -655
rect -102 -689 -86 -655
rect 86 -689 102 -655
rect 270 -689 286 -655
rect -332 -739 -298 -723
rect -332 -1131 -298 -1115
rect -74 -739 -40 -723
rect -74 -1131 -40 -1115
rect 40 -739 74 -723
rect 40 -1131 74 -1115
rect 298 -739 332 -723
rect 298 -1131 332 -1115
rect -286 -1199 -270 -1165
rect -102 -1199 -86 -1165
rect 86 -1199 102 -1165
rect 270 -1199 286 -1165
<< viali >>
rect -270 1165 -102 1199
rect 102 1165 270 1199
rect -332 795 -298 1059
rect -74 739 -40 1115
rect 40 739 74 1115
rect 298 795 332 1059
rect -270 655 -102 689
rect 102 655 270 689
rect -270 547 -102 581
rect 102 547 270 581
rect -332 177 -298 441
rect -74 121 -40 497
rect 40 121 74 497
rect 298 177 332 441
rect -270 37 -102 71
rect 102 37 270 71
rect -270 -71 -102 -37
rect 102 -71 270 -37
rect -332 -441 -298 -177
rect -74 -497 -40 -121
rect 40 -497 74 -121
rect 298 -441 332 -177
rect -270 -581 -102 -547
rect 102 -581 270 -547
rect -270 -689 -102 -655
rect 102 -689 270 -655
rect -332 -1059 -298 -795
rect -74 -1115 -40 -739
rect 40 -1115 74 -739
rect 298 -1059 332 -795
rect -270 -1199 -102 -1165
rect 102 -1199 270 -1165
<< metal1 >>
rect -282 1199 -90 1205
rect -282 1165 -270 1199
rect -102 1165 -90 1199
rect -282 1159 -90 1165
rect 90 1199 282 1205
rect 90 1165 102 1199
rect 270 1165 282 1199
rect 90 1159 282 1165
rect -80 1115 -34 1127
rect -338 1059 -292 1071
rect -338 795 -332 1059
rect -298 795 -292 1059
rect -338 783 -292 795
rect -80 739 -74 1115
rect -40 739 -34 1115
rect -80 727 -34 739
rect 34 1115 80 1127
rect 34 739 40 1115
rect 74 739 80 1115
rect 292 1059 338 1071
rect 292 795 298 1059
rect 332 795 338 1059
rect 292 783 338 795
rect 34 727 80 739
rect -282 689 -90 695
rect -282 655 -270 689
rect -102 655 -90 689
rect -282 649 -90 655
rect 90 689 282 695
rect 90 655 102 689
rect 270 655 282 689
rect 90 649 282 655
rect -282 581 -90 587
rect -282 547 -270 581
rect -102 547 -90 581
rect -282 541 -90 547
rect 90 581 282 587
rect 90 547 102 581
rect 270 547 282 581
rect 90 541 282 547
rect -80 497 -34 509
rect -338 441 -292 453
rect -338 177 -332 441
rect -298 177 -292 441
rect -338 165 -292 177
rect -80 121 -74 497
rect -40 121 -34 497
rect -80 109 -34 121
rect 34 497 80 509
rect 34 121 40 497
rect 74 121 80 497
rect 292 441 338 453
rect 292 177 298 441
rect 332 177 338 441
rect 292 165 338 177
rect 34 109 80 121
rect -282 71 -90 77
rect -282 37 -270 71
rect -102 37 -90 71
rect -282 31 -90 37
rect 90 71 282 77
rect 90 37 102 71
rect 270 37 282 71
rect 90 31 282 37
rect -282 -37 -90 -31
rect -282 -71 -270 -37
rect -102 -71 -90 -37
rect -282 -77 -90 -71
rect 90 -37 282 -31
rect 90 -71 102 -37
rect 270 -71 282 -37
rect 90 -77 282 -71
rect -80 -121 -34 -109
rect -338 -177 -292 -165
rect -338 -441 -332 -177
rect -298 -441 -292 -177
rect -338 -453 -292 -441
rect -80 -497 -74 -121
rect -40 -497 -34 -121
rect -80 -509 -34 -497
rect 34 -121 80 -109
rect 34 -497 40 -121
rect 74 -497 80 -121
rect 292 -177 338 -165
rect 292 -441 298 -177
rect 332 -441 338 -177
rect 292 -453 338 -441
rect 34 -509 80 -497
rect -282 -547 -90 -541
rect -282 -581 -270 -547
rect -102 -581 -90 -547
rect -282 -587 -90 -581
rect 90 -547 282 -541
rect 90 -581 102 -547
rect 270 -581 282 -547
rect 90 -587 282 -581
rect -282 -655 -90 -649
rect -282 -689 -270 -655
rect -102 -689 -90 -655
rect -282 -695 -90 -689
rect 90 -655 282 -649
rect 90 -689 102 -655
rect 270 -689 282 -655
rect 90 -695 282 -689
rect -80 -739 -34 -727
rect -338 -795 -292 -783
rect -338 -1059 -332 -795
rect -298 -1059 -292 -795
rect -338 -1071 -292 -1059
rect -80 -1115 -74 -739
rect -40 -1115 -34 -739
rect -80 -1127 -34 -1115
rect 34 -739 80 -727
rect 34 -1115 40 -739
rect 74 -1115 80 -739
rect 292 -795 338 -783
rect 292 -1059 298 -795
rect 332 -1059 338 -795
rect 292 -1071 338 -1059
rect 34 -1127 80 -1115
rect -282 -1165 -90 -1159
rect -282 -1199 -270 -1165
rect -102 -1199 -90 -1165
rect -282 -1205 -90 -1199
rect 90 -1165 282 -1159
rect 90 -1199 102 -1165
rect 270 -1199 282 -1165
rect 90 -1205 282 -1199
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 4 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 70 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
