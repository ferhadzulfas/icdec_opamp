magic
tech sky130A
magscale 1 2
timestamp 1729245215
<< ndiff >>
rect 688 706 742 1106
rect -54 88 0 488
<< psubdiff >>
rect -288 1225 -228 1259
rect 916 1225 976 1259
rect -288 1199 -254 1225
rect 942 1199 976 1225
rect -288 -31 -254 -5
rect 942 -31 976 -5
rect -288 -65 -228 -31
rect 916 -65 976 -31
<< psubdiffcont >>
rect -228 1225 916 1259
rect -288 -5 -254 1199
rect 942 -5 976 1199
rect -228 -65 916 -31
<< poly >>
rect -142 684 -112 694
rect -204 668 -112 684
rect -204 634 -188 668
rect -154 634 -112 668
rect -204 618 -112 634
rect 800 684 830 706
rect 800 668 892 684
rect 800 634 842 668
rect 876 634 892 668
rect -204 560 -112 576
rect -204 526 -188 560
rect -154 526 -112 560
rect 58 554 630 628
rect 800 618 892 634
rect 800 560 892 576
rect -204 510 -112 526
rect -142 488 -112 510
rect 800 526 842 560
rect 876 526 892 560
rect 800 510 892 526
rect 800 502 830 510
<< polycont >>
rect -188 634 -154 668
rect 842 634 876 668
rect -188 526 -154 560
rect 842 526 876 560
<< locali >>
rect -288 1225 -228 1259
rect 916 1225 976 1259
rect -288 1199 -254 1225
rect 942 1199 976 1225
rect -204 634 -188 668
rect -154 634 -138 668
rect 826 634 842 668
rect 876 634 892 668
rect -204 526 -188 560
rect -154 526 -138 560
rect 826 526 842 560
rect 876 526 892 560
rect -288 -31 -254 -5
rect 942 -31 976 -5
rect -288 -65 -228 -31
rect 916 -65 976 -31
<< viali >>
rect 270 1225 305 1259
rect -188 634 -154 668
rect 842 634 876 668
rect -188 526 -154 560
rect 842 526 876 560
rect 384 -65 418 -31
<< metal1 >>
rect 258 1259 317 1265
rect 258 1225 270 1259
rect 305 1225 317 1259
rect 258 1219 317 1225
rect -194 706 54 1106
rect 271 1081 305 1219
rect 636 1094 882 1106
rect 365 718 375 1094
rect 427 718 437 1094
rect 636 718 688 1094
rect 742 718 882 1094
rect -188 674 -154 706
rect 5 674 52 706
rect -200 668 -142 674
rect -200 634 -188 668
rect -154 634 -142 668
rect -200 628 -142 634
rect 5 628 104 674
rect 261 627 313 718
rect 636 706 882 718
rect 842 674 876 706
rect 830 668 888 674
rect 830 634 842 668
rect 876 634 888 668
rect 830 628 888 634
rect 261 570 427 627
rect -200 560 -142 566
rect -200 526 -188 560
rect -154 526 -142 560
rect -200 520 -142 526
rect -188 490 -154 520
rect -194 476 -60 490
rect 375 476 427 570
rect 830 560 888 566
rect 601 508 683 554
rect 830 526 842 560
rect 876 526 888 560
rect 830 520 888 526
rect 635 488 683 508
rect 842 488 876 520
rect -194 100 -54 476
rect 0 100 52 476
rect -194 88 52 100
rect -112 76 52 88
rect 251 76 261 476
rect 313 76 323 476
rect 384 -25 419 110
rect 635 90 882 488
rect 635 77 793 90
rect 372 -31 430 -25
rect 372 -65 384 -31
rect 418 -65 430 -31
rect 372 -71 430 -65
<< via1 >>
rect 375 718 427 1094
rect 688 718 742 1094
rect -54 100 0 476
rect 261 76 313 476
<< metal2 >>
rect 375 1094 427 1104
rect 375 627 427 718
rect 687 1094 743 1104
rect 687 708 743 718
rect 261 575 427 627
rect -55 476 1 486
rect -55 90 1 100
rect 261 476 313 575
rect 261 66 313 76
<< via2 >>
rect 687 718 688 1094
rect 688 718 742 1094
rect 742 718 743 1094
rect -55 100 -54 476
rect -54 100 0 476
rect 0 100 1 476
<< metal3 >>
rect 677 1094 753 1099
rect 677 718 687 1094
rect 743 718 753 1094
rect 677 628 753 718
rect -65 568 753 628
rect -65 476 11 568
rect 628 567 753 568
rect -65 100 -55 476
rect 1 100 11 476
rect -65 95 11 100
use sky130_fd_pr__nfet_01v8_6C7GGL  sky130_fd_pr__nfet_01v8_6C7GGL_0
timestamp 1729223951
transform 1 0 -127 0 1 906
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_6C7GGL  sky130_fd_pr__nfet_01v8_6C7GGL_1
timestamp 1729223951
transform 1 0 815 0 1 288
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_6C7GGL  sky130_fd_pr__nfet_01v8_6C7GGL_2
timestamp 1729223951
transform 1 0 815 0 1 906
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_6C7GGL  sky130_fd_pr__nfet_01v8_6C7GGL_3
timestamp 1729223951
transform 1 0 -127 0 1 288
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_46AA6M  sky130_fd_pr__nfet_01v8_46AA6M_0
timestamp 1729223494
transform 1 0 344 0 1 597
box -344 -597 344 597
<< labels >>
flabel metal1 282 1151 284 1154 0 FreeSans 640 0 0 0 GND
port 0 nsew
flabel metal1 30 657 32 660 0 FreeSans 640 0 0 0 D3
port 1 nsew
flabel metal2 391 666 393 669 0 FreeSans 640 0 0 0 RS
port 2 nsew
flabel metal3 701 650 703 653 0 FreeSans 640 0 0 0 D4
port 3 nsew
<< end >>
