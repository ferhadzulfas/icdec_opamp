magic
tech sky130A
magscale 1 2
timestamp 1729382277
<< psubdiff >>
rect -214 525 -154 559
rect 1435 525 1495 559
rect -214 499 -180 525
rect 1461 499 1495 525
rect -214 -610 -180 -584
rect 1461 -610 1495 -584
rect -214 -644 -154 -610
rect 1435 -644 1495 -610
<< psubdiffcont >>
rect -154 525 1435 559
rect -214 -584 -180 499
rect 1461 -584 1495 499
rect -154 -644 1435 -610
<< poly >>
rect -37 79 -7 100
rect -99 63 -7 79
rect -99 29 -83 63
rect -49 29 -7 63
rect -99 13 -7 29
rect 1265 79 1295 93
rect 1265 63 1358 79
rect 1265 29 1308 63
rect 1342 29 1358 63
rect 1265 13 1358 29
rect -99 -96 -7 -81
rect -99 -130 -83 -96
rect -49 -130 -7 -96
rect -99 -146 -7 -130
rect -37 -148 -7 -146
rect 1265 -97 1357 -81
rect 1265 -131 1307 -97
rect 1341 -131 1357 -97
rect 1265 -147 1357 -131
rect 1265 -149 1295 -147
<< polycont >>
rect -83 29 -49 63
rect 1308 29 1342 63
rect -83 -130 -49 -96
rect 1307 -131 1341 -97
<< locali >>
rect -214 525 -154 559
rect 1435 525 1495 559
rect -214 499 -180 525
rect 1461 499 1495 525
rect -99 29 -83 63
rect -49 29 -33 63
rect 1292 29 1308 63
rect 1342 29 1358 63
rect -99 -130 -83 -96
rect -49 -130 -33 -96
rect 1291 -131 1307 -97
rect 1341 -131 1357 -97
rect -214 -610 -180 -584
rect 1461 -610 1495 -584
rect -214 -644 -154 -610
rect 1435 -644 1495 -610
<< viali >>
rect -83 29 -49 63
rect 1308 29 1342 63
rect -83 -130 -49 -96
rect 1307 -131 1341 -97
rect 270 -610 325 -609
rect 270 -644 325 -610
rect 933 -644 988 -610
rect 933 -645 988 -644
<< metal1 >>
rect 591 451 601 456
rect -43 409 601 451
rect -43 301 -1 409
rect 591 404 601 409
rect 657 451 667 456
rect 657 409 1300 451
rect 657 404 667 409
rect 1258 301 1300 409
rect -89 101 45 301
rect 217 101 377 301
rect 549 101 709 301
rect 881 101 1041 301
rect 1213 101 1347 301
rect -83 69 -49 101
rect -95 63 -37 69
rect -95 29 -83 63
rect -49 29 -37 63
rect -95 23 -37 29
rect 70 20 80 72
rect 182 20 192 72
rect -95 -96 -37 -90
rect -95 -130 -83 -96
rect -49 -130 -37 -96
rect -95 -136 -37 -130
rect -83 -171 -49 -136
rect 70 -140 80 -88
rect 182 -140 192 -88
rect 269 -168 325 101
rect 600 73 659 101
rect 593 72 603 73
rect 402 69 524 72
rect 592 69 603 72
rect 400 23 603 69
rect 402 20 524 23
rect 592 20 603 23
rect 593 19 603 20
rect 657 69 667 73
rect 734 69 856 72
rect 657 23 858 69
rect 657 19 667 23
rect 734 20 856 23
rect 402 -140 412 -88
rect 514 -140 524 -88
rect 734 -140 744 -88
rect 846 -140 856 -88
rect 933 -168 989 101
rect 1066 20 1076 72
rect 1178 20 1188 72
rect 1307 69 1342 101
rect 1296 63 1354 69
rect 1296 29 1308 63
rect 1342 29 1354 63
rect 1296 23 1354 29
rect 1066 -140 1076 -88
rect 1178 -140 1188 -88
rect 1295 -97 1353 -91
rect 1295 -131 1307 -97
rect 1341 -131 1353 -97
rect 1295 -137 1353 -131
rect -82 -180 -49 -171
rect -43 -181 -1 -169
rect -58 -357 -48 -181
rect 4 -357 14 -181
rect -43 -477 -1 -357
rect 217 -368 269 -168
rect 259 -369 269 -368
rect 325 -368 377 -168
rect 591 -169 601 -168
rect 325 -369 335 -368
rect 549 -369 601 -169
rect 657 -169 667 -168
rect 923 -169 933 -168
rect 657 -369 709 -169
rect 881 -369 933 -169
rect 989 -169 999 -168
rect 1307 -169 1341 -137
rect 989 -369 1041 -169
rect 1213 -181 1347 -169
rect 1213 -357 1254 -181
rect 1306 -357 1347 -181
rect 1213 -369 1347 -357
rect 1259 -477 1301 -369
rect -43 -519 1301 -477
rect 260 -603 270 -600
rect 258 -650 270 -603
rect 325 -603 335 -600
rect 260 -652 270 -650
rect 325 -650 337 -603
rect 923 -604 933 -601
rect 325 -652 335 -650
rect 921 -651 933 -604
rect 988 -604 998 -601
rect 923 -653 933 -651
rect 988 -651 1000 -604
rect 988 -653 998 -651
<< via1 >>
rect 601 404 657 456
rect 80 20 182 72
rect 80 -140 182 -88
rect 603 19 657 73
rect 412 -140 514 -88
rect 744 -140 846 -88
rect 1076 20 1178 72
rect 1076 -140 1178 -88
rect -48 -357 4 -181
rect 269 -369 325 -168
rect 601 -369 657 -168
rect 933 -369 989 -168
rect 1254 -357 1306 -181
rect 270 -609 325 -600
rect 270 -644 325 -609
rect 270 -652 325 -644
rect 933 -610 988 -601
rect 933 -645 988 -610
rect 933 -653 988 -645
<< metal2 >>
rect 601 458 657 468
rect 601 392 657 402
rect 80 72 182 82
rect 80 -30 182 20
rect 603 73 657 83
rect 1076 72 1178 82
rect 657 19 658 25
rect 603 -30 658 19
rect 1076 -30 1178 20
rect -48 -88 1306 -30
rect -48 -181 4 -88
rect 80 -150 182 -140
rect 412 -150 514 -140
rect 744 -150 846 -140
rect 1076 -150 1178 -140
rect -48 -367 4 -357
rect 269 -168 325 -158
rect 269 -379 325 -369
rect 601 -168 657 -158
rect 601 -379 657 -369
rect 933 -168 989 -158
rect 1254 -181 1306 -88
rect 1254 -367 1306 -357
rect 933 -379 989 -369
rect 270 -469 325 -379
rect 933 -469 988 -379
rect 270 -524 988 -469
rect 270 -600 325 -524
rect 270 -662 325 -652
rect 933 -601 988 -524
rect 933 -663 988 -653
<< via2 >>
rect 601 456 657 458
rect 601 404 657 456
rect 601 402 657 404
rect 601 -369 657 -168
<< metal3 >>
rect 591 458 667 463
rect 591 402 601 458
rect 657 402 667 458
rect 591 -168 667 402
rect 591 -369 601 -168
rect 657 -369 667 -168
rect 591 -374 667 -369
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1729382277
transform 1 0 1280 0 1 -269
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1729382277
transform 1 0 -22 0 1 -269
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1729382277
transform 1 0 -22 0 1 201
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1729382277
transform 1 0 1280 0 1 201
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_H42E3S  sky130_fd_pr__nfet_01v8_H42E3S_0
timestamp 1729324418
transform 1 0 629 0 1 -269
box -636 -188 636 188
use sky130_fd_pr__nfet_01v8_H42E3S  sky130_fd_pr__nfet_01v8_H42E3S_1
timestamp 1729324418
transform 1 0 629 0 1 201
box -636 -188 636 188
<< labels >>
flabel metal2 140 -56 140 -56 0 FreeSans 640 0 0 0 D6
port 0 nsew
flabel metal3 623 -134 623 -134 0 FreeSans 640 0 0 0 OUT
port 1 nsew
flabel metal2 967 -562 967 -562 0 FreeSans 640 0 0 0 GND
port 2 nsew
<< end >>
