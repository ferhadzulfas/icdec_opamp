magic
tech sky130A
magscale 1 2
timestamp 1729236971
<< error_p >>
rect -36 399 36 405
rect -36 365 -24 399
rect -36 359 36 365
rect -144 18 144 236
rect -36 -37 36 -31
rect -36 -71 -24 -37
rect -36 -77 36 -71
rect -36 -365 36 -359
rect -36 -399 -24 -365
rect -36 -405 36 -399
<< nwell >>
rect -144 18 144 418
rect -144 -418 144 -18
<< pmos >>
rect -50 118 50 318
rect -50 -318 50 -118
<< pdiff >>
rect -108 306 -50 318
rect -108 130 -96 306
rect -62 130 -50 306
rect -108 118 -50 130
rect 50 306 108 318
rect 50 130 62 306
rect 96 130 108 306
rect 50 118 108 130
rect -108 -130 -50 -118
rect -108 -306 -96 -130
rect -62 -306 -50 -130
rect -108 -318 -50 -306
rect 50 -130 108 -118
rect 50 -306 62 -130
rect 96 -306 108 -130
rect 50 -318 108 -306
<< pdiffc >>
rect -96 130 -62 306
rect 62 130 96 306
rect -96 -306 -62 -130
rect 62 -306 96 -130
<< poly >>
rect -50 399 50 415
rect -50 365 -34 399
rect 34 365 50 399
rect -50 318 50 365
rect -50 71 50 118
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -118 50 -71
rect -50 -365 50 -318
rect -50 -399 -34 -365
rect 34 -399 50 -365
rect -50 -415 50 -399
<< polycont >>
rect -34 365 34 399
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -399 34 -365
<< locali >>
rect -50 365 -34 399
rect 34 365 50 399
rect -96 306 -62 322
rect -96 114 -62 130
rect 62 306 96 322
rect 62 114 96 130
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -130 -62 -114
rect -96 -322 -62 -306
rect 62 -130 96 -114
rect 62 -322 96 -306
rect -50 -399 -34 -365
rect 34 -399 50 -365
<< viali >>
rect -24 365 24 399
rect -96 130 -62 306
rect 62 130 96 306
rect -24 37 24 71
rect -24 -71 24 -37
rect -96 -306 -62 -130
rect 62 -306 96 -130
rect -24 -399 24 -365
<< metal1 >>
rect -36 399 36 405
rect -36 365 -24 399
rect 24 365 36 399
rect -36 359 36 365
rect -102 306 -56 318
rect -102 130 -96 306
rect -62 130 -56 306
rect -102 118 -56 130
rect 56 306 102 318
rect 56 130 62 306
rect 96 130 102 306
rect 56 118 102 130
rect -36 71 36 77
rect -36 37 -24 71
rect 24 37 36 71
rect -36 31 36 37
rect -36 -37 36 -31
rect -36 -71 -24 -37
rect 24 -71 36 -37
rect -36 -77 36 -71
rect -102 -130 -56 -118
rect -102 -306 -96 -130
rect -62 -306 -56 -130
rect -102 -318 -56 -306
rect 56 -130 102 -118
rect 56 -306 62 -130
rect 96 -306 102 -130
rect 56 -318 102 -306
rect -36 -365 36 -359
rect -36 -399 -24 -365
rect 24 -399 36 -365
rect -36 -405 36 -399
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 2 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
