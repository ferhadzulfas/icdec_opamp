magic
tech sky130A
magscale 1 2
timestamp 1729324418
<< nmos >>
rect -578 -100 -418 100
rect -246 -100 -86 100
rect 86 -100 246 100
rect 418 -100 578 100
<< ndiff >>
rect -636 88 -578 100
rect -636 -88 -624 88
rect -590 -88 -578 88
rect -636 -100 -578 -88
rect -418 88 -360 100
rect -418 -88 -406 88
rect -372 -88 -360 88
rect -418 -100 -360 -88
rect -304 88 -246 100
rect -304 -88 -292 88
rect -258 -88 -246 88
rect -304 -100 -246 -88
rect -86 88 -28 100
rect -86 -88 -74 88
rect -40 -88 -28 88
rect -86 -100 -28 -88
rect 28 88 86 100
rect 28 -88 40 88
rect 74 -88 86 88
rect 28 -100 86 -88
rect 246 88 304 100
rect 246 -88 258 88
rect 292 -88 304 88
rect 246 -100 304 -88
rect 360 88 418 100
rect 360 -88 372 88
rect 406 -88 418 88
rect 360 -100 418 -88
rect 578 88 636 100
rect 578 -88 590 88
rect 624 -88 636 88
rect 578 -100 636 -88
<< ndiffc >>
rect -624 -88 -590 88
rect -406 -88 -372 88
rect -292 -88 -258 88
rect -74 -88 -40 88
rect 40 -88 74 88
rect 258 -88 292 88
rect 372 -88 406 88
rect 590 -88 624 88
<< poly >>
rect -578 172 -418 188
rect -578 138 -562 172
rect -434 138 -418 172
rect -578 100 -418 138
rect -246 172 -86 188
rect -246 138 -230 172
rect -102 138 -86 172
rect -246 100 -86 138
rect 86 172 246 188
rect 86 138 102 172
rect 230 138 246 172
rect 86 100 246 138
rect 418 172 578 188
rect 418 138 434 172
rect 562 138 578 172
rect 418 100 578 138
rect -578 -138 -418 -100
rect -578 -172 -562 -138
rect -434 -172 -418 -138
rect -578 -188 -418 -172
rect -246 -138 -86 -100
rect -246 -172 -230 -138
rect -102 -172 -86 -138
rect -246 -188 -86 -172
rect 86 -138 246 -100
rect 86 -172 102 -138
rect 230 -172 246 -138
rect 86 -188 246 -172
rect 418 -138 578 -100
rect 418 -172 434 -138
rect 562 -172 578 -138
rect 418 -188 578 -172
<< polycont >>
rect -562 138 -434 172
rect -230 138 -102 172
rect 102 138 230 172
rect 434 138 562 172
rect -562 -172 -434 -138
rect -230 -172 -102 -138
rect 102 -172 230 -138
rect 434 -172 562 -138
<< locali >>
rect -578 138 -562 172
rect -434 138 -418 172
rect -246 138 -230 172
rect -102 138 -86 172
rect 86 138 102 172
rect 230 138 246 172
rect 418 138 434 172
rect 562 138 578 172
rect -624 88 -590 104
rect -624 -104 -590 -88
rect -406 88 -372 104
rect -406 -104 -372 -88
rect -292 88 -258 104
rect -292 -104 -258 -88
rect -74 88 -40 104
rect -74 -104 -40 -88
rect 40 88 74 104
rect 40 -104 74 -88
rect 258 88 292 104
rect 258 -104 292 -88
rect 372 88 406 104
rect 372 -104 406 -88
rect 590 88 624 104
rect 590 -104 624 -88
rect -578 -172 -562 -138
rect -434 -172 -418 -138
rect -246 -172 -230 -138
rect -102 -172 -86 -138
rect 86 -172 102 -138
rect 230 -172 246 -138
rect 418 -172 434 -138
rect 562 -172 578 -138
<< viali >>
rect -549 138 -447 172
rect -217 138 -115 172
rect 115 138 217 172
rect 447 138 549 172
rect -624 -88 -590 88
rect -406 -88 -372 88
rect -292 -88 -258 88
rect -74 -88 -40 88
rect 40 -88 74 88
rect 258 -88 292 88
rect 372 -88 406 88
rect 590 -88 624 88
rect -549 -172 -447 -138
rect -217 -172 -115 -138
rect 115 -172 217 -138
rect 447 -172 549 -138
<< metal1 >>
rect -561 172 -435 178
rect -561 138 -549 172
rect -447 138 -435 172
rect -561 132 -435 138
rect -229 172 -103 178
rect -229 138 -217 172
rect -115 138 -103 172
rect -229 132 -103 138
rect 103 172 229 178
rect 103 138 115 172
rect 217 138 229 172
rect 103 132 229 138
rect 435 172 561 178
rect 435 138 447 172
rect 549 138 561 172
rect 435 132 561 138
rect -630 88 -584 100
rect -630 -88 -624 88
rect -590 -88 -584 88
rect -630 -100 -584 -88
rect -412 88 -366 100
rect -412 -88 -406 88
rect -372 -88 -366 88
rect -412 -100 -366 -88
rect -298 88 -252 100
rect -298 -88 -292 88
rect -258 -88 -252 88
rect -298 -100 -252 -88
rect -80 88 -34 100
rect -80 -88 -74 88
rect -40 -88 -34 88
rect -80 -100 -34 -88
rect 34 88 80 100
rect 34 -88 40 88
rect 74 -88 80 88
rect 34 -100 80 -88
rect 252 88 298 100
rect 252 -88 258 88
rect 292 -88 298 88
rect 252 -100 298 -88
rect 366 88 412 100
rect 366 -88 372 88
rect 406 -88 412 88
rect 366 -100 412 -88
rect 584 88 630 100
rect 584 -88 590 88
rect 624 -88 630 88
rect 584 -100 630 -88
rect -561 -138 -435 -132
rect -561 -172 -549 -138
rect -447 -172 -435 -138
rect -561 -178 -435 -172
rect -229 -138 -103 -132
rect -229 -172 -217 -138
rect -115 -172 -103 -138
rect -229 -178 -103 -172
rect 103 -138 229 -132
rect 103 -172 115 -138
rect 217 -172 229 -138
rect 103 -178 229 -172
rect 435 -138 561 -132
rect 435 -172 447 -138
rect 549 -172 561 -138
rect 435 -178 561 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
