magic
tech sky130A
magscale 1 2
timestamp 1729387919
<< nwell >>
rect 94 -2032 894 512
<< nsubdiff >>
rect 131 442 226 476
rect 765 442 858 476
rect 131 399 165 442
rect 824 399 858 442
rect 131 -1962 165 -1919
rect 824 -1962 858 -1919
rect 131 -1996 226 -1962
rect 765 -1996 858 -1962
<< nsubdiffcont >>
rect 226 442 765 476
rect 131 -1919 165 399
rect 824 -1919 858 399
rect 226 -1996 765 -1962
<< poly >>
rect 278 -150 308 -109
rect 216 -166 308 -150
rect 216 -200 232 -166
rect 266 -200 308 -166
rect 216 -216 308 -200
rect 682 -149 712 -118
rect 682 -165 774 -149
rect 682 -199 724 -165
rect 758 -199 774 -165
rect 682 -215 774 -199
rect 278 -644 308 -603
rect 216 -660 308 -644
rect 216 -694 232 -660
rect 266 -694 308 -660
rect 216 -710 308 -694
rect 682 -643 712 -601
rect 682 -659 774 -643
rect 682 -693 724 -659
rect 758 -693 774 -659
rect 216 -806 308 -790
rect 216 -840 232 -806
rect 266 -840 308 -806
rect 366 -809 466 -699
rect 524 -809 624 -699
rect 682 -709 774 -693
rect 682 -805 773 -789
rect 216 -856 308 -840
rect 278 -884 308 -856
rect 682 -839 723 -805
rect 757 -839 773 -805
rect 682 -855 773 -839
rect 682 -890 712 -855
rect 216 -1299 308 -1283
rect 216 -1333 232 -1299
rect 266 -1333 308 -1299
rect 216 -1349 308 -1333
rect 278 -1386 308 -1349
rect 682 -1299 773 -1283
rect 682 -1333 723 -1299
rect 757 -1333 773 -1299
rect 682 -1349 773 -1333
rect 682 -1382 712 -1349
<< polycont >>
rect 232 -200 266 -166
rect 724 -199 758 -165
rect 232 -694 266 -660
rect 724 -693 758 -659
rect 232 -840 266 -806
rect 723 -839 757 -805
rect 232 -1333 266 -1299
rect 723 -1333 757 -1299
<< locali >>
rect 131 442 226 476
rect 765 442 858 476
rect 131 399 165 442
rect 824 399 858 442
rect 216 -200 232 -166
rect 266 -200 282 -166
rect 708 -199 724 -165
rect 758 -199 774 -165
rect 216 -694 232 -660
rect 266 -694 282 -660
rect 708 -693 724 -659
rect 758 -693 774 -659
rect 216 -840 232 -806
rect 266 -840 282 -806
rect 707 -839 723 -805
rect 757 -839 773 -805
rect 216 -1333 232 -1299
rect 266 -1333 282 -1299
rect 707 -1333 723 -1299
rect 757 -1333 773 -1299
rect 131 -1962 165 -1919
rect 824 -1962 858 -1919
rect 131 -1996 226 -1962
rect 765 -1996 858 -1962
<< viali >>
rect 353 442 549 476
rect 232 -200 266 -166
rect 724 -199 758 -165
rect 232 -694 266 -660
rect 724 -693 758 -659
rect 232 -840 266 -806
rect 723 -839 757 -805
rect 232 -1333 266 -1299
rect 723 -1333 757 -1299
<< metal1 >>
rect 341 476 561 482
rect 341 442 353 476
rect 549 442 561 476
rect 341 436 561 442
rect 278 352 715 408
rect 774 352 784 407
rect 278 82 320 352
rect 226 -118 360 82
rect 457 -106 467 70
rect 523 -106 533 70
rect 661 -106 671 70
rect 723 -102 733 70
rect 723 -106 758 -102
rect 232 -160 266 -118
rect 220 -166 278 -160
rect 220 -200 232 -166
rect 266 -200 278 -166
rect 220 -206 278 -200
rect 382 -236 450 -198
rect 530 -208 540 -156
rect 608 -208 618 -156
rect 724 -159 758 -106
rect 712 -165 770 -159
rect 712 -199 724 -165
rect 758 -199 770 -165
rect 712 -205 770 -199
rect 382 -289 608 -236
rect 372 -374 382 -322
rect 450 -374 460 -322
rect 540 -332 608 -289
rect 226 -424 360 -413
rect 630 -424 764 -412
rect 213 -600 223 -424
rect 275 -600 360 -424
rect 457 -600 467 -424
rect 523 -600 533 -424
rect 630 -600 715 -424
rect 767 -600 777 -424
rect 226 -612 360 -600
rect 630 -612 764 -600
rect 232 -654 266 -612
rect 724 -653 758 -612
rect 220 -660 278 -654
rect 220 -694 232 -660
rect 266 -694 278 -660
rect 220 -700 278 -694
rect 712 -659 770 -653
rect 712 -693 724 -659
rect 758 -693 770 -659
rect 712 -699 770 -693
rect 220 -806 278 -800
rect 220 -840 232 -806
rect 266 -840 278 -806
rect 220 -846 278 -840
rect 711 -805 769 -799
rect 711 -839 723 -805
rect 757 -839 769 -805
rect 711 -845 769 -839
rect 232 -906 266 -846
rect 723 -906 758 -845
rect 226 -918 360 -906
rect 630 -918 764 -906
rect 213 -1094 223 -918
rect 275 -1094 360 -918
rect 460 -1094 470 -918
rect 522 -1094 532 -918
rect 630 -1094 715 -918
rect 767 -1094 777 -918
rect 226 -1106 360 -1094
rect 630 -1106 764 -1094
rect 372 -1196 382 -1144
rect 450 -1196 460 -1144
rect 540 -1224 608 -1185
rect 383 -1243 608 -1224
rect 382 -1272 608 -1243
rect 220 -1299 278 -1293
rect 220 -1333 232 -1299
rect 266 -1333 278 -1299
rect 382 -1319 450 -1272
rect 711 -1299 769 -1293
rect 220 -1339 278 -1333
rect 232 -1400 266 -1339
rect 530 -1362 540 -1310
rect 608 -1362 618 -1310
rect 711 -1333 723 -1299
rect 757 -1333 769 -1299
rect 711 -1339 769 -1333
rect 226 -1600 360 -1400
rect 459 -1588 469 -1412
rect 521 -1588 531 -1412
rect 661 -1588 671 -1412
rect 723 -1416 758 -1339
rect 723 -1588 733 -1416
rect 278 -1875 330 -1600
rect 278 -1931 715 -1875
rect 771 -1931 781 -1875
<< via1 >>
rect 715 352 774 407
rect 467 -106 523 70
rect 671 -106 723 70
rect 540 -208 608 -156
rect 382 -374 450 -322
rect 223 -600 275 -424
rect 467 -600 523 -424
rect 715 -600 767 -424
rect 223 -1094 275 -918
rect 470 -1094 522 -918
rect 715 -1094 767 -918
rect 382 -1196 450 -1144
rect 540 -1362 608 -1310
rect 469 -1588 521 -1412
rect 671 -1588 723 -1412
rect 715 -1931 771 -1875
<< metal2 >>
rect 716 417 772 418
rect 715 408 774 417
rect 715 407 716 408
rect 772 407 774 408
rect 715 342 774 352
rect 215 248 713 306
rect 215 109 279 248
rect 216 -424 278 109
rect 671 80 713 248
rect 467 70 523 80
rect 467 -116 523 -106
rect 671 70 723 80
rect 671 -116 723 -106
rect 540 -156 608 -146
rect 540 -232 608 -208
rect 382 -282 608 -232
rect 382 -322 450 -282
rect 382 -384 450 -374
rect 216 -600 223 -424
rect 275 -600 278 -424
rect 216 -918 278 -600
rect 467 -424 523 -414
rect 467 -610 523 -600
rect 713 -424 769 -414
rect 713 -610 769 -600
rect 216 -1094 223 -918
rect 275 -1094 278 -918
rect 216 -1765 278 -1094
rect 467 -918 523 -908
rect 467 -1104 523 -1094
rect 715 -918 771 -908
rect 715 -1104 771 -1094
rect 382 -1144 450 -1134
rect 382 -1220 450 -1196
rect 382 -1269 608 -1220
rect 540 -1310 608 -1269
rect 540 -1372 608 -1362
rect 467 -1412 523 -1402
rect 467 -1598 523 -1588
rect 671 -1412 723 -1402
rect 671 -1598 723 -1588
rect 671 -1765 712 -1598
rect 216 -1826 712 -1765
rect 715 -1875 771 -1865
rect 715 -1941 771 -1931
<< via2 >>
rect 716 407 772 408
rect 716 352 772 407
rect 467 -106 523 70
rect 467 -600 523 -424
rect 713 -600 715 -424
rect 715 -600 767 -424
rect 767 -600 769 -424
rect 467 -1094 470 -918
rect 470 -1094 522 -918
rect 522 -1094 523 -918
rect 715 -1094 767 -918
rect 767 -1094 771 -918
rect 467 -1588 469 -1412
rect 469 -1588 521 -1412
rect 521 -1588 523 -1412
rect 715 -1931 771 -1875
<< metal3 >>
rect 706 408 782 413
rect 706 352 716 408
rect 772 352 782 408
rect 706 347 782 352
rect 457 70 533 75
rect 457 -106 467 70
rect 523 -106 533 70
rect 457 -111 533 -106
rect 465 -419 525 -111
rect 712 -419 774 347
rect 457 -424 533 -419
rect 457 -600 467 -424
rect 523 -600 533 -424
rect 457 -605 533 -600
rect 703 -424 779 -419
rect 703 -600 713 -424
rect 769 -600 779 -424
rect 703 -605 779 -600
rect 465 -913 525 -605
rect 712 -913 774 -605
rect 457 -918 533 -913
rect 457 -1094 467 -918
rect 523 -1094 533 -918
rect 457 -1099 533 -1094
rect 705 -918 781 -913
rect 705 -1094 715 -918
rect 771 -1094 781 -918
rect 705 -1099 781 -1094
rect 465 -1407 525 -1099
rect 457 -1412 533 -1407
rect 457 -1588 467 -1412
rect 523 -1588 533 -1412
rect 712 -1588 774 -1099
rect 457 -1593 533 -1588
rect 713 -1870 774 -1588
rect 705 -1875 781 -1870
rect 705 -1931 715 -1875
rect 771 -1931 781 -1875
rect 705 -1936 781 -1931
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729236971
transform 1 0 293 0 1 -1500
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729236971
transform 1 0 697 0 1 -18
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729236971
transform 1 0 293 0 1 -18
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1729236971
transform 1 0 293 0 1 -512
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729236971
transform 1 0 697 0 1 -512
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729236971
transform 1 0 293 0 1 -1006
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729236971
transform 1 0 697 0 1 -1006
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_8
timestamp 1729236971
transform 1 0 697 0 1 -1500
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_VQXXLL  sky130_fd_pr__pfet_01v8_VQXXLL_0
timestamp 1729236971
transform 1 0 495 0 1 -18
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXXLL  sky130_fd_pr__pfet_01v8_VQXXLL_1
timestamp 1729236971
transform 1 0 495 0 1 -512
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXXLL  sky130_fd_pr__pfet_01v8_VQXXLL_2
timestamp 1729236971
transform 1 0 495 0 1 -1006
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXXLL  sky130_fd_pr__pfet_01v8_VQXXLL_3
timestamp 1729236971
transform 1 0 495 0 1 -1500
box -223 -200 223 200
<< labels >>
flabel viali 476 464 476 464 0 FreeSans 640 0 0 0 VDD
port 0 nsew
flabel metal1 416 368 416 368 0 FreeSans 640 0 0 0 OUT
port 1 nsew
flabel metal2 472 278 472 278 0 FreeSans 640 0 0 0 D6
port 2 nsew
flabel metal1 404 -218 404 -218 0 FreeSans 640 0 0 0 VIP
port 3 nsew
flabel metal2 422 -302 422 -302 0 FreeSans 640 0 0 0 VIN
port 4 nsew
flabel metal3 494 -398 494 -398 0 FreeSans 640 0 0 0 D5
port 6 nsew
<< end >>
